////////////////////////////////////////////////////////////////////////////////
// Company     : XnonymouX
//
// Filename    : mux2
// Description : 2:1 parallel mux.
//
// Author      : Duong Nguyen
// Created On  : 10-6-2015
// History     : Initial 	
//
////////////////////////////////////////////////////////////////////////////////

module mux2
    (
    //-------------------
    //In 0
    sel0,
    in0,
    //-------------------
    //In 1
    sel1,
    in1,
    //-------------------
    //Out
    out
    );

//------------------------------------------------------------------------------
//Parameters
parameter DW = 1'b1;
//------------------------------------------------------------------------------
// Port declarations
input               sel0;
input [DW-1:0]	    in0;
//
input               sel1;
input [DW-1:0]	    in1;
//
output [DW-1:0]	    out;
//------------------------------------------------------------------------------
//internal signal

//------------------------------------------------------------------------------
//Logic
assign out = ({DW{sel0}} & in0) |
             ({DW{sel1}} & in1);

endmodule 

