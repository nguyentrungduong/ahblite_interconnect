////////////////////////////////////////////////////////////////////////////////
// Company     : XnonymouX
//
// Filename    : mux9
// Description : 9:1 parallel mux.
//
// Author      : Duong Nguyen
// Created On  : 10-6-2015
// History     : Initial 	
//
////////////////////////////////////////////////////////////////////////////////

module mux9
    (
    sel0,
    in0,
    //-------------------
    sel1,
    in1,
    //-------------------
    sel2,
    in2,
    //-------------------
    sel3,
    in3,
    //-------------------
    sel4,
    in4,
    //-------------------
    sel5,
    in5,
    //-------------------
    sel6,
    in6,
    //-------------------
    sel7,
    in7,
    //-------------------
    sel8,
    in8,
    //-------------------
    out
    );

//------------------------------------------------------------------------------
//Parameters
parameter DW = 1'b1;
//------------------------------------------------------------------------------
// Port declarations
input               sel0;
input [DW-1:0]	    in0;
//
input               sel1;
input [DW-1:0]	    in1;
//
input               sel2;
input [DW-1:0]	    in2;
//
input               sel3;
input [DW-1:0]	    in3;
//
input               sel4;
input [DW-1:0]	    in4;
//
input               sel5;
input [DW-1:0]	    in5;
//
input               sel6;
input [DW-1:0]	    in6;
//
input               sel7;
input [DW-1:0]	    in7;
//
input               sel8;
input [DW-1:0]	    in8;
//
output [DW-1:0]	    out;
//------------------------------------------------------------------------------
//internal signal
wire [DW-1:0]       out04;
wire [DW-1:0]       out58;
//------------------------------------------------------------------------------
//Mux 5:1
mux5   #(.DW(DW))   mux5_0 
    (
    .sel0  (sel0),
    .in0   (in0),
    //-------------------
    .sel1  (sel1),
    .in1   (in1),
    //-------------------
    .sel2  (sel2),
    .in2   (in2),
    //-------------------
    .sel3  (sel3),
    .in3   (in3),
    //-------------------
    .sel4  (sel4),
    .in4   (in4),
    //-------------------
    .out   (out04)
    );
//------------------------------------------------------------------------------
//Mux 4:1
mux4   #(.DW(DW))   mux4_0 
    (
    .sel0  (sel5),
    .in0   (in5),
    //-------------------
    .sel1  (sel6),
    .in1   (in6),
    //-------------------
    .sel2  (sel7),
    .in2   (in7),
    //-------------------
    .sel3  (sel8),
    .in3   (in8),
    //-------------------
    .out   (out58)
    );
//------------------------------------------------------------------------------
//Mux 2:1
assign out = out04 | out58;

endmodule 

